`timescale 1ns / 100ps
/**
 * 
 * Todo:
 *  - MUX for the end-points;
 *  - MUX-select for the end-points;
 */
module enc_datapath
  ( input clock,
    input reset,

    input s1_tvalid,
    input s2_tvalid,
    input s3_tvalid,
    input s4_tvalid
    );


endmodule  /* enc_datapath */
