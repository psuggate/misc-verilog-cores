`timescale 1ns / 100ps
module ddr3_top_tb;

endmodule  // ddr3_top_tb
